package serialalu_pkg;
	import uvm_pkg::*;

	`include "serialalu_sequencer.sv"
	`include "serialalu_monitor.sv"
	`include "serialalu_driver.sv"
	`include "serialalu_agent.sv"
	`include "serialalu_scoreboard.sv"
	`include "serialalu_config.sv"
	`include "serialalu_env.sv"
	`include "serialalu_test.sv"
endpackage: serialalu_pkg
